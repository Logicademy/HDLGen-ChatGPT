-- Header Section
-- Component Name : test
-- Title          : 
-- Description    : 
-- Author(s)      : 
-- Company        : 
-- Email          : 
-- Date           : 13/07/2022


-- Library Section
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

