-- Package
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
package MainPackage is
type array4x32 is array(3 downto 0) of std_logic_vector(31 downto 0);
type array5x32 is array(4 downto 0) of signed(31 downto 0);
type array6x32 is array(5 downto 0) of unsigned(31 downto 0);


end MainPackage;
package body MainPackage is
end MainPackage;

