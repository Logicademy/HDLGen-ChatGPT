// Note on arrays in Verilog
//
// <FM> if verilog and HDLGen defines an array port signal, e.g, [m:n] XYZ [p:q]
// Assume q = 0 and n = 0
// r = p+1, o = m+1, ro = r*0
// merge the signal as [ro-1:0] XYZ_'r*o' in module

// Example
// <FM> Here [31:0] reg4x32_CSRA [3:0], m=31, n=0, p=3, q=0, r=4, o=32, ro=128
// merge the signal as [127:0] reg4x32_CSRA_128 in module
// Define input  input  [127:0] reg4x32_CSRA_128;
// Define internal array signal 
// wire [31:0] reg4x32_CSRA [3:0];
// In testbench, use the 128 bit signal
// If the component is used in a hierarchical design, can assign an array in the next level (to the merged vector) and process in the next level as an array




/* 
   Header section
   Generated by HDLGen, Github https://github.com/abishek-bupathi/HDLGen
   Reference: https://tinyurl.com/VerilogTips 
      
   Component Name : threshold
   Title          : Generate a 32-x32-bit threshold array from 32x32-byte source data array
*/

/*
   Description
   Generate a 32-x32-bit threshold array from 
   - 32x32-byte source data array
   - threshVal(7:0)

   Result bit is asserted if souce byte >= threshVal

   Author(s)      : Fearghal Morgan
   Company        : University of Galway
   Email          : fearghal.morgan@universityofgalway.ie
   Date           : 29/03/2023
*/

/*
   module signal dictionary
   clk  System clock strobe
   rst  Asynchronous reset signal, asserted h 
   ce	threshold component enable. Assertion (h) activates the threshold register components.
   go	Assertion (h) activates threshold finite state machine (FSM)
   reg4x32_CSRA	4 x 32-bit register memory, control and status register A
   reg4x32_CSRB	4 x 32-bit register memory, control and status register B
   BRAM_dOut	256-bit block RAM (BRAM) memory
   active	Asserted to highlight that FSM is active. Signal is a flag and is not used externally. 
   wr	Assertion (h) synchronously writes memory(add) = dataToMem(31:0)
   add	memory address
   datToMem	memory write data
   functBus	96-bit bus which can be connected to any threshold component signals, to be stored / viewed during threshold function execution
*/

/* 
  internal signal dictionary
   NS 	Finite State Machine (FSM) next state and current state
   CS 	Finite State Machine (FSM) next state and current state 
   NSYAdd	Y address std_logic_vector state signals
   CSYAdd	Y address std_logic_vector state signals
   NSXAdd	X address std_logic_vector state signals
   CSXAdd	X address std_logic_vector state signals
   BRAMByte	BRAM_dOut(CSXAdd*8+7 : CSXAdd*8)
   NSThreshVec	thresholdVec std_logic_vector state signals
   CSThreshVec	thresholdVec std_logic_vector state signals
   threshVal	threshVal(7:0) = reg4x32_CSRA(31:24)
*/

// FM No library declarations required //

// module declaration
module threshold(
		clk,
		rst,
		ce,
		go,
		reg4x32_CSRA_128,
		reg4x32_CSRB_128,
		BRAM_dOut,
		
		active,
		wr,
		add,
		datToMem,
		functBus
	);

// <FM> outdent port definitions to left margin
// Port definitions
input  clk;
input  rst;
input  ce;
input  go;
input  [127:0] reg4x32_CSRA_128;
input  [127:0] reg4x32_CSRB_128;
input  [255:0] BRAM_dOut;

output active;
output wr;
output [7:0] add;
output [31:0] datToMem;
output [95:0] functBus;

// Internal signal declarations
// Use localparam approach since it is more compact
//   parameter idle = 2'b00;
//   parameter chkBRAM_Byte_GT_thresholdValue = 2'b01;
//   parameter wr_threshVec_to_reg32x32 = 2'b10;
//   parameter write_status_to_reg4x32_CSRA0 = 2'b11;

// Internal signal declarations

// Declare states 
localparam [1:0]
idle = 0, 
chkBRAM_Byte_GT_thresholdValue = 1, 
wr_threshVec_to_reg32x32 = 2, 
write_status_to_reg4x32_CSRA0 = 3;
	
reg active;
reg wr;
reg [7:0] add;
reg [31:0] datToMem;

reg [1:0] NS;
reg [1:0] CS;    
reg [4:0]  NSYAdd;
reg [4:0]  CSYAdd;
reg [4:0]  NSXAdd;
reg [4:0]  CSXAdd;
reg [31:0] NSThreshVec;
reg [31:0] CSThreshVec;
wire [7:0]  BRAMByte;
wire [7:0]  threshVal;

// handling arrays: create internal array signal
wire [31:0] reg4x32_CSRA [3:0]; 
wire [31:0] reg4x32_CSRB [3:0]; 
 
// FM automate generation of array from concatentation port vector signal
// assign {reg4x32_CSRA[3],reg4x32_CSRA[2],reg4x32_CSRA[1],reg4x32_CSRA[0]} = reg4x32_CSRA_128;
assign reg4x32_CSRA[3] = reg4x32_CSRA_128[127:96];
assign reg4x32_CSRA[2] = reg4x32_CSRA_128[95:64];
assign reg4x32_CSRA[1] = reg4x32_CSRA_128[63:32];
assign reg4x32_CSRA[0] = reg4x32_CSRA_128[31:0];
// assign {reg4x32_CSRB[3],reg4x32_CSRB[2],reg4x32_CSRB[1],reg4x32_CSRB[0]} = reg4x32_CSRB_128;
assign reg4x32_CSRB[3] = reg4x32_CSRB_128[127:96];
assign reg4x32_CSRB[2] = reg4x32_CSRB_128[95:64];
assign reg4x32_CSRB[1] = reg4x32_CSRB_128[63:32];
assign reg4x32_CSRB[0] = reg4x32_CSRB_128[31:0];
 
// Assign internal signals
assign BRAMByte = BRAM_dOut[CSXAdd*8 +:8];// take 8 bit slice, starting at bit CSXAdd*8
assign threshVal = reg4x32_CSRA[0][15:8]; // check indices 
	
// Assign output signals
assign functBus = 128'h0;
    
    // stateReg 
    always @(posedge clk or posedge rst) 
     begin : stateReg
    	// Complete the process if required
    	if ( rst ) 
		 begin
    		CS <= idle;
    		CSYAdd <= 5'b0;
    		CSXAdd <= 5'b0;
    		CSThreshVec <= 32'b0;
    	 end
		else
		 begin
		    if (ce)
    	 	 begin 
    		  CS <= NS;
    		  CSYAdd <= NSYAdd;
    		  CSXAdd <= NSXAdd;
    		  CSThreshVec <= NSThreshVec;
    		 end
	     end 
     end
    
    // NSAndOPDecode 
    // Complete the process if required
	always @(CS or go or reg4x32_CSRA[0] or reg4x32_CSRB[0] or CSYAdd or CSXAdd or CSThreshVec or threshVal or BRAMByte)
   	  begin : NSAndOPDecode
        NS     <= CS;   // default
        active <= 1'b1; // default asserted
        NSYAdd <= CSYAdd;
        NSXAdd <= CSXAdd;
        NSThreshVec <= CSThreshVec;
        wr <= 1'b0; 
        add <= {3'b010, CSYAdd}; // address 32 x 256-bit BRAM
	    datToMem <= CSThreshVec;

    	case ( CS )
    		idle:
    			begin
     		      NSYAdd <= 0; 
    		      NSXAdd <= 0;
    		      NSThreshVec <= 0; 
				  // assign other output signal states
                  if (go) 
                    begin
                      NS <= chkBRAM_Byte_GT_thresholdValue;
					  add <= {3'b010, CSYAdd}; // address 32 x 256-bit BRAM
                    end
				  else
				    begin
	      		      active <= 1'b0;
					end
    			end

    		 chkBRAM_Byte_GT_thresholdValue:
    			begin 
				  add <= {3'b010, CSYAdd}; // address 32 x 256-bit BRAM
			      if (BRAMByte > threshVal)      
			        begin
			          NSThreshVec[CSXAdd] <= 1'b1; // set single bit of vector
			        end 
			      NSXAdd <= CSXAdd + 1;   // increment XAdd counter
				  if (NSXAdd == 31)
				    begin
				      NS <= wr_threshVec_to_reg32x32; // final threshVec value is ready in wr_threshVec_to_reg32x32 state
				    end 
				end

    		 wr_threshVec_to_reg32x32:
    			begin
    		      wr <= 1'b1; 
                  add <= {3'b001, CSYAdd}; // resultMem address
                  datToMem <= CSThreshVec;
                  NS <= write_status_to_reg4x32_CSRA0;
	              NSThreshVec <= 0;
			      NSYAdd <= CSYAdd + 1;        // increment YAdd counter
		          NS <= chkBRAM_Byte_GT_thresholdValue; // loop, to process next BRAM word
	   		      if (NSYAdd == 31) 
				    NS <= write_status_to_reg4x32_CSRA0;    // final threshVec value is ready in wr_threshVec_to_reg32x32 state
    			 end

    		 write_status_to_reg4x32_CSRA0:
    			begin
    		      wr <= 1'b1; 
				  add <= 8'b0; // address CSRA[0]
                  datToMem <= {reg4x32_CSRA[0][31:2], 2'b10};
                  NS <= idle;
    			end
								
    		default:
    			begin
    			end
    	endcase
      end

endmodule