-- Header Section
-- Component Name : mux21_1
-- Title          : To be Completedkhlerjkllkerj

-- Description
-- To be Completedoed
-- dhildclkh

-- Author(s)      : jp
-- Company        : ug
-- Email          : lkhlklk
-- Date           : 04/10/2022

-- entity signal dictionary
-- select	jkrlkj
-- jkfeckjl	to be completed

-- internal signal dictionary
-- None

-- library declarations
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

-- entity declaration
entity mux21_1 is 
Port(
	select : in std_logic;
	jkfeckjl : out std_logic
);
end entity mux21_1;

architecture Combinational of mux21_1 is
-- Internal signal declarations

-- Component declarations

begin

jkrfj: process(select)
begin
	-- Complete the process
	jkfeckjl <= select;

end process;

end Combinational;