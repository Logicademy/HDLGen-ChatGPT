-- Package
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
package arrayPackage is


end arrayPackage;
package body arrayPackage is
end arrayPackage;

